magic
tech sky130A
timestamp 1702697407
<< nwell >>
rect -135 770 635 910
<< nmos >>
rect 0 535 30 635
rect 80 535 110 635
rect 160 535 175 635
rect 225 535 255 635
rect 305 535 335 635
rect 385 535 400 635
rect 450 535 480 635
rect 530 535 560 635
rect 0 0 15 100
rect 65 0 80 100
rect 130 0 145 100
rect 195 0 210 100
rect 260 0 275 100
rect 325 0 340 100
rect 390 0 420 100
rect 470 0 500 100
rect 550 0 565 100
<< pmos >>
rect -65 790 -50 890
rect 80 790 95 890
rect 120 790 135 890
rect 185 790 200 890
rect 445 790 460 890
rect 510 790 525 890
rect 550 790 565 890
<< ndiff >>
rect -50 620 0 635
rect -50 550 -35 620
rect -15 550 0 620
rect -50 535 0 550
rect 30 620 80 635
rect 30 550 45 620
rect 65 550 80 620
rect 30 535 80 550
rect 110 620 160 635
rect 110 550 125 620
rect 145 550 160 620
rect 110 535 160 550
rect 175 620 225 635
rect 175 550 190 620
rect 210 550 225 620
rect 175 535 225 550
rect 255 620 305 635
rect 255 550 270 620
rect 290 550 305 620
rect 255 535 305 550
rect 335 620 385 635
rect 335 550 350 620
rect 370 550 385 620
rect 335 535 385 550
rect 400 620 450 635
rect 400 550 415 620
rect 435 550 450 620
rect 400 535 450 550
rect 480 620 530 635
rect 480 550 495 620
rect 515 550 530 620
rect 480 535 530 550
rect 560 620 610 635
rect 560 550 575 620
rect 595 550 610 620
rect 560 535 610 550
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 145 85 195 100
rect 145 15 160 85
rect 180 15 195 85
rect 145 0 195 15
rect 210 85 260 100
rect 210 15 225 85
rect 245 15 260 85
rect 210 0 260 15
rect 275 85 325 100
rect 275 15 290 85
rect 310 15 325 85
rect 275 0 325 15
rect 340 85 390 100
rect 340 15 355 85
rect 375 15 390 85
rect 340 0 390 15
rect 420 85 470 100
rect 420 15 435 85
rect 455 15 470 85
rect 420 0 470 15
rect 500 85 550 100
rect 500 15 515 85
rect 535 15 550 85
rect 500 0 550 15
rect 565 85 615 100
rect 565 15 580 85
rect 600 15 615 85
rect 565 0 615 15
<< pdiff >>
rect -115 875 -65 890
rect -115 805 -100 875
rect -80 805 -65 875
rect -115 790 -65 805
rect -50 875 0 890
rect -50 805 -35 875
rect -15 805 0 875
rect -50 790 0 805
rect 30 875 80 890
rect 30 805 45 875
rect 65 805 80 875
rect 30 790 80 805
rect 95 790 120 890
rect 135 875 185 890
rect 135 805 150 875
rect 170 805 185 875
rect 135 790 185 805
rect 200 875 250 890
rect 200 805 215 875
rect 235 805 250 875
rect 200 790 250 805
rect 395 875 445 890
rect 395 805 410 875
rect 430 805 445 875
rect 395 790 445 805
rect 460 875 510 890
rect 460 805 475 875
rect 495 805 510 875
rect 460 790 510 805
rect 525 790 550 890
rect 565 875 615 890
rect 565 805 580 875
rect 600 805 615 875
rect 565 790 615 805
<< ndiffc >>
rect -35 550 -15 620
rect 45 550 65 620
rect 125 550 145 620
rect 190 550 210 620
rect 270 550 290 620
rect 350 550 370 620
rect 415 550 435 620
rect 495 550 515 620
rect 575 550 595 620
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
rect 160 15 180 85
rect 225 15 245 85
rect 290 15 310 85
rect 355 15 375 85
rect 435 15 455 85
rect 515 15 535 85
rect 580 15 600 85
<< pdiffc >>
rect -100 805 -80 875
rect -35 805 -15 875
rect 45 805 65 875
rect 150 805 170 875
rect 215 805 235 875
rect 410 805 430 875
rect 475 805 495 875
rect 580 805 600 875
<< psubdiff >>
rect 270 705 370 720
rect 270 680 285 705
rect 355 680 370 705
rect 270 665 370 680
<< nsubdiff >>
rect 280 875 365 890
rect 280 805 295 875
rect 350 805 365 875
rect 280 790 365 805
<< psubdiffcont >>
rect 285 680 355 705
<< nsubdiffcont >>
rect 295 805 350 875
<< poly >>
rect 55 935 565 945
rect 55 915 65 935
rect 85 930 565 935
rect 85 915 95 930
rect 55 905 95 915
rect -65 890 -50 905
rect 80 890 95 905
rect 120 890 135 905
rect 185 890 200 905
rect 445 890 460 905
rect 510 890 525 905
rect 550 890 565 930
rect -65 775 -50 790
rect 80 775 95 790
rect 120 775 135 790
rect 185 775 200 790
rect 445 775 460 790
rect 510 775 525 790
rect 550 775 565 790
rect 120 765 245 775
rect 120 760 215 765
rect 205 745 215 760
rect 235 745 245 765
rect 205 735 245 745
rect 400 765 525 775
rect 400 745 410 765
rect 430 760 525 765
rect 430 745 440 760
rect 400 735 440 745
rect 0 635 30 650
rect 80 635 110 650
rect 160 635 175 650
rect 225 635 255 650
rect 305 635 335 650
rect 385 635 400 650
rect 450 635 480 650
rect 530 635 560 650
rect 0 375 30 535
rect 80 375 110 535
rect 160 480 175 535
rect 135 470 175 480
rect 135 450 145 470
rect 165 450 175 470
rect 135 440 175 450
rect 225 375 255 535
rect 305 375 335 535
rect 385 440 400 535
rect 360 430 400 440
rect 360 410 370 430
rect 390 410 400 430
rect 360 400 400 410
rect 450 375 480 535
rect 530 375 560 535
rect 0 360 560 375
rect 460 325 500 335
rect 460 305 470 325
rect 490 305 500 325
rect 460 295 500 305
rect 0 285 210 295
rect 0 265 10 285
rect 30 280 210 285
rect 30 265 40 280
rect 0 255 40 265
rect 0 100 15 255
rect 105 225 145 235
rect 105 205 115 225
rect 135 205 145 225
rect 105 195 145 205
rect 65 100 80 115
rect 130 100 145 195
rect 195 100 210 280
rect 260 185 300 195
rect 260 165 270 185
rect 290 165 300 185
rect 260 155 300 165
rect 260 100 275 155
rect 325 145 365 155
rect 325 125 335 145
rect 355 125 365 145
rect 470 125 500 295
rect 325 115 365 125
rect 325 100 340 115
rect 390 110 500 125
rect 390 100 420 110
rect 470 100 500 110
rect 550 100 565 115
rect 0 -15 15 0
rect 65 -40 80 0
rect 130 -15 145 0
rect 195 -15 210 0
rect 260 -15 275 0
rect 325 -15 340 0
rect 390 -15 420 0
rect 470 -15 500 0
rect 550 -40 565 0
rect -45 -50 565 -40
rect -45 -70 -35 -50
rect -15 -55 565 -50
rect -15 -70 -5 -55
rect -45 -80 -5 -70
<< polycont >>
rect 65 915 85 935
rect 215 745 235 765
rect 410 745 430 765
rect 145 450 165 470
rect 370 410 390 430
rect 470 305 490 325
rect 10 265 30 285
rect 115 205 135 225
rect 270 165 290 185
rect 335 125 355 145
rect -35 -70 -15 -50
<< locali >>
rect -115 935 95 945
rect -115 925 65 935
rect 55 915 65 925
rect 85 915 95 935
rect 55 905 95 915
rect -110 875 -70 885
rect -110 805 -100 875
rect -80 805 -70 875
rect -110 795 -70 805
rect -45 875 -5 885
rect -45 805 -35 875
rect -15 805 -5 875
rect -45 760 -5 805
rect -45 740 -35 760
rect -15 740 -5 760
rect -45 730 -5 740
rect 35 875 75 885
rect 35 805 45 875
rect 65 805 75 875
rect 35 760 75 805
rect 140 875 180 885
rect 140 805 150 875
rect 170 805 180 875
rect 140 795 180 805
rect 205 875 245 885
rect 205 805 215 875
rect 235 805 245 875
rect 35 740 45 760
rect 65 740 75 760
rect 35 730 75 740
rect 205 765 245 805
rect 285 875 360 885
rect 285 805 295 875
rect 350 805 360 875
rect 285 795 360 805
rect 400 875 440 885
rect 400 805 410 875
rect 430 805 440 875
rect 205 745 215 765
rect 235 745 245 765
rect 205 735 245 745
rect 400 765 440 805
rect 465 875 505 885
rect 465 805 475 875
rect 495 805 505 875
rect 465 795 505 805
rect 570 875 610 885
rect 570 805 580 875
rect 600 805 610 875
rect 400 745 410 765
rect 430 745 440 765
rect 400 735 440 745
rect 570 760 610 805
rect 570 740 580 760
rect 600 740 610 760
rect 570 730 610 740
rect 275 705 365 715
rect 275 680 285 705
rect 355 680 365 705
rect 275 670 365 680
rect -45 620 -5 630
rect -45 550 -35 620
rect -15 550 -5 620
rect -45 520 -5 550
rect 35 620 75 630
rect 35 550 45 620
rect 65 550 75 620
rect 35 540 75 550
rect 115 620 155 630
rect 115 550 125 620
rect 145 550 155 620
rect 115 520 155 550
rect -45 500 155 520
rect 180 620 220 630
rect 180 550 190 620
rect 210 550 220 620
rect 180 520 220 550
rect 260 620 300 630
rect 260 550 270 620
rect 290 550 300 620
rect 260 540 300 550
rect 340 620 380 630
rect 340 550 350 620
rect 370 550 380 620
rect 340 520 380 550
rect 180 500 380 520
rect 405 620 445 630
rect 405 550 415 620
rect 435 550 445 620
rect 405 520 445 550
rect 485 620 525 630
rect 485 550 495 620
rect 515 550 525 620
rect 485 540 525 550
rect 565 620 605 630
rect 565 550 575 620
rect 595 550 605 620
rect 565 520 605 550
rect 405 500 605 520
rect 135 470 175 480
rect 135 450 145 470
rect 165 450 175 470
rect 135 440 175 450
rect 360 430 400 440
rect 360 410 370 430
rect 390 410 400 430
rect 360 400 400 410
rect -60 325 500 335
rect -60 315 470 325
rect 460 305 470 315
rect 490 305 500 325
rect 460 295 500 305
rect -60 285 40 295
rect -60 265 10 285
rect 30 265 40 285
rect -60 255 40 265
rect -60 225 145 235
rect -60 215 115 225
rect 105 205 115 215
rect 135 205 145 225
rect 105 195 145 205
rect 260 185 465 195
rect 260 165 270 185
rect 290 175 465 185
rect 290 165 300 175
rect -45 150 -5 160
rect -45 130 -35 150
rect -15 130 -5 150
rect -45 85 -5 130
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 -50 -5 15
rect 20 150 75 160
rect 260 155 300 165
rect 20 130 45 150
rect 65 130 75 150
rect 325 145 365 155
rect 325 135 335 145
rect 20 120 75 130
rect 150 125 335 135
rect 355 125 365 145
rect 20 85 60 120
rect 150 115 365 125
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect 85 -15 125 15
rect 150 85 190 115
rect 150 15 160 85
rect 180 15 190 85
rect 150 5 190 15
rect 215 85 255 95
rect 215 15 225 85
rect 245 15 255 85
rect 215 -15 255 15
rect 280 85 320 95
rect 280 15 290 85
rect 310 15 320 85
rect 280 5 320 15
rect 345 85 385 95
rect 345 15 355 85
rect 375 15 385 85
rect 85 -35 255 -15
rect 345 -15 385 15
rect 425 85 465 175
rect 570 150 610 160
rect 570 130 580 150
rect 600 130 610 150
rect 425 15 435 85
rect 455 15 465 85
rect 425 5 465 15
rect 505 85 545 95
rect 505 15 515 85
rect 535 15 545 85
rect 505 -15 545 15
rect 570 85 610 130
rect 570 15 580 85
rect 600 15 610 85
rect 570 5 610 15
rect 345 -35 545 -15
rect -45 -70 -35 -50
rect -15 -70 -5 -50
rect -45 -80 -5 -70
<< viali >>
rect -100 805 -80 875
rect -35 740 -15 760
rect 150 805 170 875
rect 45 740 65 760
rect 295 805 350 875
rect 475 805 495 875
rect 580 740 600 760
rect 45 550 65 620
rect 270 550 290 620
rect 495 550 515 620
rect -35 130 -15 150
rect 45 130 65 150
rect 290 15 310 85
rect 580 130 600 150
<< metal1 >>
rect -115 875 615 890
rect -115 805 -100 875
rect -80 805 150 875
rect 170 805 295 875
rect 350 805 475 875
rect 495 805 615 875
rect -115 790 615 805
rect -50 770 0 775
rect -50 730 -45 770
rect -5 730 0 770
rect -50 635 0 730
rect 30 770 80 775
rect 30 730 35 770
rect 75 730 80 770
rect 30 635 80 730
rect 565 770 615 775
rect 565 730 570 770
rect 610 730 615 770
rect 270 635 370 720
rect 565 635 615 730
rect -50 620 615 635
rect -50 550 45 620
rect 65 550 270 620
rect 290 550 495 620
rect 515 550 615 620
rect -50 535 615 550
rect -50 160 0 535
rect -50 120 -45 160
rect -5 120 0 160
rect -50 115 0 120
rect 30 160 80 535
rect 30 120 35 160
rect 75 120 80 160
rect 30 115 80 120
rect 565 160 615 535
rect 565 120 570 160
rect 610 120 615 160
rect 565 115 615 120
rect -50 85 615 100
rect -50 15 290 85
rect 310 15 615 85
rect -50 0 615 15
<< via1 >>
rect -45 760 -5 770
rect -45 740 -35 760
rect -35 740 -15 760
rect -15 740 -5 760
rect -45 730 -5 740
rect 35 760 75 770
rect 35 740 45 760
rect 45 740 65 760
rect 65 740 75 760
rect 35 730 75 740
rect 570 760 610 770
rect 570 740 580 760
rect 580 740 600 760
rect 600 740 610 760
rect 570 730 610 740
rect -45 150 -5 160
rect -45 130 -35 150
rect -35 130 -15 150
rect -15 130 -5 150
rect -45 120 -5 130
rect 35 150 75 160
rect 35 130 45 150
rect 45 130 65 150
rect 65 130 75 150
rect 35 120 75 130
rect 570 150 610 160
rect 570 130 580 150
rect 580 130 600 150
rect 600 130 610 150
rect 570 120 610 130
<< metal2 >>
rect -50 770 0 775
rect -50 730 -45 770
rect -5 730 0 770
rect -50 160 0 730
rect -50 120 -45 160
rect -5 120 0 160
rect -50 115 0 120
rect 30 770 80 775
rect 30 730 35 770
rect 75 730 80 770
rect 30 160 80 730
rect 30 120 35 160
rect 75 120 80 160
rect 30 115 80 120
rect 565 770 615 775
rect 565 730 570 770
rect 610 730 615 770
rect 565 160 615 730
rect 565 120 570 160
rect 610 120 615 160
rect 565 115 615 120
<< end >>
