magic
tech sky130A
timestamp 1702528739
<< nwell >>
rect -130 225 380 365
rect 275 220 380 225
rect 275 20 365 220
<< nmos >>
rect -60 45 -45 145
rect 5 45 20 145
rect 170 45 185 145
rect -60 -180 -45 -80
rect 5 -180 20 -80
rect 45 -180 60 -80
rect 110 -180 125 -80
rect 150 -180 165 -80
rect 215 -180 230 -80
<< pmos >>
rect -60 245 -45 345
rect 5 245 20 345
rect 45 245 60 345
rect 190 245 205 345
rect 230 245 245 345
rect 295 245 310 345
<< ndiff >>
rect -110 130 -60 145
rect -110 60 -95 130
rect -75 60 -60 130
rect -110 45 -60 60
rect -45 130 5 145
rect -45 60 -30 130
rect -10 60 5 130
rect -45 45 5 60
rect 20 130 70 145
rect 120 130 170 145
rect 20 60 35 130
rect 55 60 70 130
rect 120 60 135 130
rect 155 60 170 130
rect 20 45 70 60
rect 120 45 170 60
rect 185 130 235 145
rect 185 60 200 130
rect 220 60 235 130
rect 185 45 235 60
rect -110 -95 -60 -80
rect -110 -165 -95 -95
rect -75 -165 -60 -95
rect -110 -180 -60 -165
rect -45 -95 5 -80
rect -45 -165 -30 -95
rect -10 -165 5 -95
rect -45 -180 5 -165
rect 20 -180 45 -80
rect 60 -95 110 -80
rect 60 -165 75 -95
rect 95 -165 110 -95
rect 60 -180 110 -165
rect 125 -180 150 -80
rect 165 -95 215 -80
rect 165 -165 180 -95
rect 200 -165 215 -95
rect 165 -180 215 -165
rect 230 -95 280 -80
rect 230 -165 245 -95
rect 265 -165 280 -95
rect 230 -180 280 -165
<< pdiff >>
rect -110 330 -60 345
rect -110 260 -95 330
rect -75 260 -60 330
rect -110 245 -60 260
rect -45 330 5 345
rect -45 260 -30 330
rect -10 260 5 330
rect -45 245 5 260
rect 20 245 45 345
rect 60 330 110 345
rect 60 260 75 330
rect 95 260 110 330
rect 60 245 110 260
rect 140 330 190 345
rect 140 260 155 330
rect 175 260 190 330
rect 140 245 190 260
rect 205 245 230 345
rect 245 330 295 345
rect 245 260 260 330
rect 280 260 295 330
rect 245 245 295 260
rect 310 330 360 345
rect 310 260 325 330
rect 345 260 360 330
rect 310 245 360 260
<< ndiffc >>
rect -95 60 -75 130
rect -30 60 -10 130
rect 35 60 55 130
rect 135 60 155 130
rect 200 60 220 130
rect -95 -165 -75 -95
rect -30 -165 -10 -95
rect 75 -165 95 -95
rect 180 -165 200 -95
rect 245 -165 265 -95
<< pdiffc >>
rect -95 260 -75 330
rect -30 260 -10 330
rect 75 260 95 330
rect 155 260 175 330
rect 260 260 280 330
rect 325 260 345 330
<< psubdiff >>
rect 70 130 120 145
rect 70 60 90 130
rect 110 60 120 130
rect 70 45 120 60
<< nsubdiff >>
rect 295 130 345 145
rect 295 60 310 130
rect 330 60 345 130
rect 295 45 345 60
<< psubdiffcont >>
rect 90 60 110 130
<< nsubdiffcont >>
rect 310 60 330 130
<< poly >>
rect 95 390 135 395
rect 95 370 105 390
rect 125 370 135 390
rect -60 345 -45 360
rect 5 345 20 360
rect 45 355 205 370
rect 45 345 60 355
rect 190 345 205 355
rect 230 345 245 360
rect 295 345 310 360
rect -60 235 -45 245
rect 5 235 20 245
rect -60 225 20 235
rect 45 230 60 245
rect 190 230 205 245
rect 230 235 245 245
rect 295 235 310 245
rect -85 220 20 225
rect 230 220 310 235
rect -85 200 -75 220
rect -55 200 -45 220
rect -85 195 -45 200
rect 270 200 280 220
rect 300 200 310 220
rect 270 195 310 200
rect -110 155 -45 170
rect -60 145 -45 155
rect 5 145 20 160
rect 170 145 185 160
rect -60 30 -45 45
rect 5 30 20 45
rect 170 30 185 45
rect -115 20 -85 30
rect -115 0 -110 20
rect -90 5 -85 20
rect -90 0 230 5
rect -115 -10 230 0
rect -85 -40 -45 -35
rect -85 -60 -75 -40
rect -55 -60 -45 -40
rect -85 -65 -45 -60
rect -60 -80 -45 -65
rect 5 -80 20 -65
rect 45 -80 60 -65
rect 110 -80 125 -65
rect 150 -80 165 -65
rect 215 -80 230 -10
rect -60 -195 -45 -180
rect 5 -245 20 -180
rect 45 -190 60 -180
rect 110 -190 125 -180
rect 45 -200 125 -190
rect 45 -205 75 -200
rect 65 -220 75 -205
rect 95 -205 125 -200
rect 95 -220 105 -205
rect 65 -225 105 -220
rect -20 -250 20 -245
rect -20 -270 -10 -250
rect 10 -270 20 -250
rect -20 -275 20 -270
rect 150 -245 165 -180
rect 215 -195 230 -180
rect 150 -250 190 -245
rect 150 -270 160 -250
rect 180 -270 190 -250
rect 150 -275 190 -270
<< polycont >>
rect 105 370 125 390
rect -75 200 -55 220
rect 280 200 300 220
rect -110 0 -90 20
rect -75 -60 -55 -40
rect 75 -220 95 -200
rect -10 -270 10 -250
rect 160 -270 180 -250
<< locali >>
rect 95 390 135 395
rect -130 370 105 390
rect 125 370 135 390
rect 95 365 135 370
rect -105 330 -65 340
rect -105 260 -95 330
rect -75 260 -65 330
rect -105 250 -65 260
rect -40 330 0 340
rect -40 260 -30 330
rect -10 260 0 330
rect -40 250 0 260
rect 65 330 105 340
rect 65 260 75 330
rect 95 260 105 330
rect 65 250 105 260
rect 145 330 185 340
rect 145 260 155 330
rect 175 260 185 330
rect 145 250 185 260
rect 250 330 290 340
rect 250 260 260 330
rect 280 260 290 330
rect 250 250 290 260
rect 315 330 355 340
rect 315 260 325 330
rect 345 260 355 330
rect 315 250 355 260
rect -95 225 -75 250
rect -95 220 -45 225
rect -95 200 -75 220
rect -55 200 -45 220
rect -95 195 -45 200
rect 270 220 310 225
rect 270 200 280 220
rect 300 200 310 220
rect 270 195 310 200
rect -95 145 -75 195
rect 270 180 290 195
rect 35 160 290 180
rect -105 130 -65 145
rect 35 140 55 160
rect -105 60 -95 130
rect -75 60 -65 130
rect -105 50 -65 60
rect -40 130 0 140
rect -40 60 -30 130
rect -10 60 0 130
rect -40 50 0 60
rect 25 130 65 140
rect 25 60 35 130
rect 55 60 65 130
rect 25 50 65 60
rect 85 130 165 140
rect 85 60 90 130
rect 110 60 135 130
rect 155 60 165 130
rect 85 50 165 60
rect 190 130 230 140
rect 190 60 200 130
rect 220 60 230 130
rect 190 50 230 60
rect 300 130 340 140
rect 300 60 310 130
rect 330 60 340 130
rect 300 50 340 60
rect -30 30 -10 50
rect 200 30 220 50
rect -115 20 -85 30
rect -115 0 -110 20
rect -90 0 -85 20
rect -30 10 220 30
rect -115 -10 -85 0
rect -25 -25 5 -15
rect -115 -40 -45 -35
rect -115 -60 -75 -40
rect -55 -60 -45 -40
rect -25 -45 -20 -25
rect 0 -45 5 -25
rect -25 -55 5 -45
rect -115 -65 -45 -60
rect -105 -95 -65 -85
rect -105 -165 -95 -95
rect -75 -165 -65 -95
rect -105 -195 -65 -165
rect -40 -95 0 -85
rect -40 -165 -30 -95
rect -10 -165 0 -95
rect -40 -175 0 -165
rect 65 -95 105 -85
rect 65 -165 75 -95
rect 95 -165 105 -95
rect 65 -175 105 -165
rect 170 -95 210 -85
rect 170 -165 180 -95
rect 200 -165 210 -95
rect 170 -175 210 -165
rect 235 -95 275 -85
rect 235 -165 245 -95
rect 265 -165 275 -95
rect 235 -195 275 -165
rect -105 -200 275 -195
rect -105 -220 75 -200
rect 95 -220 275 -200
rect -105 -225 275 -220
rect -130 -250 290 -245
rect -130 -270 -10 -250
rect 10 -270 160 -250
rect 180 -270 290 -250
rect -130 -275 290 -270
<< viali >>
rect -30 260 -10 330
rect 260 260 280 330
rect 90 60 110 130
rect 135 60 155 130
rect 310 60 330 130
rect -20 -45 0 -25
rect 75 -165 95 -95
<< metal1 >>
rect -130 330 380 340
rect -130 260 -30 330
rect -10 260 260 330
rect 280 260 380 330
rect -130 250 380 260
rect 85 130 165 140
rect 85 60 90 130
rect 110 60 135 130
rect 155 60 165 130
rect 85 50 165 60
rect 300 130 340 140
rect 300 60 310 130
rect 330 60 340 130
rect 300 50 340 60
rect -25 -25 5 -15
rect -25 -45 -20 -25
rect 0 -45 5 -25
rect -25 -55 5 -45
rect -130 -95 285 -85
rect -130 -165 75 -95
rect 95 -165 285 -95
rect -130 -175 285 -165
<< end >>
