magic
tech sky130A
timestamp 1702700917
<< nwell >>
rect -135 735 635 875
<< nmos >>
rect 0 535 30 635
rect 80 535 110 635
rect 160 535 175 635
rect 225 535 255 635
rect 305 535 335 635
rect 385 535 400 635
rect 450 535 480 635
rect 530 535 560 635
rect 0 0 15 100
rect 65 0 80 100
rect 130 0 145 100
rect 195 0 210 100
rect 260 0 275 100
rect 325 0 340 100
rect 390 0 420 100
rect 470 0 500 100
rect 550 0 565 100
<< pmos >>
rect -65 755 -50 855
rect 80 755 95 855
rect 120 755 135 855
rect 185 755 200 855
rect 445 755 460 855
rect 510 755 525 855
rect 550 755 565 855
<< ndiff >>
rect -50 620 0 635
rect -50 550 -35 620
rect -15 550 0 620
rect -50 535 0 550
rect 30 620 80 635
rect 30 550 45 620
rect 65 550 80 620
rect 30 535 80 550
rect 110 620 160 635
rect 110 550 125 620
rect 145 550 160 620
rect 110 535 160 550
rect 175 620 225 635
rect 175 550 190 620
rect 210 550 225 620
rect 175 535 225 550
rect 255 620 305 635
rect 255 550 270 620
rect 290 550 305 620
rect 255 535 305 550
rect 335 620 385 635
rect 335 550 350 620
rect 370 550 385 620
rect 335 535 385 550
rect 400 620 450 635
rect 400 550 415 620
rect 435 550 450 620
rect 400 535 450 550
rect 480 620 530 635
rect 480 550 495 620
rect 515 550 530 620
rect 480 535 530 550
rect 560 620 610 635
rect 560 550 575 620
rect 595 550 610 620
rect 560 535 610 550
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 145 85 195 100
rect 145 15 160 85
rect 180 15 195 85
rect 145 0 195 15
rect 210 85 260 100
rect 210 15 225 85
rect 245 15 260 85
rect 210 0 260 15
rect 275 85 325 100
rect 275 15 290 85
rect 310 15 325 85
rect 275 0 325 15
rect 340 85 390 100
rect 340 15 355 85
rect 375 15 390 85
rect 340 0 390 15
rect 420 85 470 100
rect 420 15 435 85
rect 455 15 470 85
rect 420 0 470 15
rect 500 85 550 100
rect 500 15 515 85
rect 535 15 550 85
rect 500 0 550 15
rect 565 85 615 100
rect 565 15 580 85
rect 600 15 615 85
rect 565 0 615 15
<< pdiff >>
rect -115 840 -65 855
rect -115 770 -100 840
rect -80 770 -65 840
rect -115 755 -65 770
rect -50 840 0 855
rect -50 770 -35 840
rect -15 770 0 840
rect -50 755 0 770
rect 30 840 80 855
rect 30 770 45 840
rect 65 770 80 840
rect 30 755 80 770
rect 95 755 120 855
rect 135 840 185 855
rect 135 770 150 840
rect 170 770 185 840
rect 135 755 185 770
rect 200 840 250 855
rect 200 770 215 840
rect 235 770 250 840
rect 200 755 250 770
rect 395 840 445 855
rect 395 770 410 840
rect 430 770 445 840
rect 395 755 445 770
rect 460 840 510 855
rect 460 770 475 840
rect 495 770 510 840
rect 460 755 510 770
rect 525 755 550 855
rect 565 840 615 855
rect 565 770 580 840
rect 600 770 615 840
rect 565 755 615 770
<< ndiffc >>
rect -35 550 -15 620
rect 45 550 65 620
rect 125 550 145 620
rect 190 550 210 620
rect 270 550 290 620
rect 350 550 370 620
rect 415 550 435 620
rect 495 550 515 620
rect 575 550 595 620
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
rect 160 15 180 85
rect 225 15 245 85
rect 290 15 310 85
rect 355 15 375 85
rect 435 15 455 85
rect 515 15 535 85
rect 580 15 600 85
<< pdiffc >>
rect -100 770 -80 840
rect -35 770 -15 840
rect 45 770 65 840
rect 150 770 170 840
rect 215 770 235 840
rect 410 770 430 840
rect 475 770 495 840
rect 580 770 600 840
<< psubdiff >>
rect 270 705 370 720
rect 270 680 285 705
rect 355 680 370 705
rect 270 665 370 680
<< nsubdiff >>
rect 280 840 365 855
rect 280 770 295 840
rect 350 770 365 840
rect 280 755 365 770
<< psubdiffcont >>
rect 285 680 355 705
<< nsubdiffcont >>
rect 295 770 350 840
<< poly >>
rect 55 900 565 910
rect 55 880 65 900
rect 85 895 565 900
rect 85 880 95 895
rect 55 870 95 880
rect -65 855 -50 870
rect 80 855 95 870
rect 120 855 135 870
rect 185 855 200 870
rect 445 855 460 870
rect 510 855 525 870
rect 550 855 565 895
rect -65 735 -50 755
rect 80 740 95 755
rect 120 740 135 755
rect 185 740 200 755
rect 445 740 460 755
rect 510 740 525 755
rect 550 740 565 755
rect -65 725 -5 735
rect 120 730 245 740
rect 120 725 215 730
rect -65 720 -35 725
rect -45 705 -35 720
rect -15 705 -5 725
rect -45 695 -5 705
rect 205 710 215 725
rect 235 710 245 730
rect 400 730 525 740
rect 205 700 245 710
rect 400 710 410 730
rect 430 725 525 730
rect 430 710 440 725
rect 400 700 440 710
rect 0 635 30 650
rect 80 635 110 650
rect 160 635 175 650
rect 225 635 255 650
rect 305 635 335 650
rect 385 635 400 650
rect 450 635 480 650
rect 530 635 560 650
rect 0 375 30 535
rect 80 375 110 535
rect 160 480 175 535
rect 135 470 175 480
rect 135 450 145 470
rect 165 450 175 470
rect 135 440 175 450
rect 225 375 255 535
rect 305 375 335 535
rect 385 440 400 535
rect 360 430 400 440
rect 360 410 370 430
rect 390 410 400 430
rect 360 400 400 410
rect 450 375 480 535
rect 530 400 560 535
rect 520 390 560 400
rect 520 375 530 390
rect 0 370 530 375
rect 550 370 560 390
rect 0 360 560 370
rect 460 325 500 335
rect 460 305 470 325
rect 490 305 500 325
rect 460 295 500 305
rect 0 285 210 295
rect 0 265 10 285
rect 30 280 210 285
rect 30 265 40 280
rect 0 255 40 265
rect 0 100 15 255
rect 105 225 145 235
rect 105 205 115 225
rect 135 205 145 225
rect 105 195 145 205
rect 65 100 80 115
rect 130 100 145 195
rect 195 100 210 280
rect 260 185 300 195
rect 260 165 270 185
rect 290 165 300 185
rect 260 155 300 165
rect 260 100 275 155
rect 325 145 365 155
rect 325 125 335 145
rect 355 125 365 145
rect 470 125 500 295
rect 325 115 365 125
rect 325 100 340 115
rect 390 110 500 125
rect 390 100 420 110
rect 470 100 500 110
rect 550 100 565 115
rect 0 -15 15 0
rect 65 -40 80 0
rect 130 -15 145 0
rect 195 -15 210 0
rect 260 -15 275 0
rect 325 -15 340 0
rect 390 -15 420 0
rect 470 -15 500 0
rect 550 -40 565 0
rect -45 -50 565 -40
rect -45 -70 -35 -50
rect -15 -55 565 -50
rect -15 -70 -5 -55
rect -45 -80 -5 -70
<< polycont >>
rect 65 880 85 900
rect -35 705 -15 725
rect 215 710 235 730
rect 410 710 430 730
rect 145 450 165 470
rect 370 410 390 430
rect 530 370 550 390
rect 470 305 490 325
rect 10 265 30 285
rect 115 205 135 225
rect 270 165 290 185
rect 335 125 355 145
rect -35 -70 -15 -50
<< locali >>
rect -135 900 95 910
rect -135 890 65 900
rect 55 880 65 890
rect 85 880 95 900
rect 55 870 95 880
rect -110 840 -70 850
rect -110 770 -100 840
rect -80 770 -70 840
rect -110 760 -70 770
rect -45 840 -5 850
rect -45 770 -35 840
rect -15 770 -5 840
rect -45 725 -5 770
rect -45 705 -35 725
rect -15 705 -5 725
rect -45 695 -5 705
rect 35 840 75 850
rect 35 770 45 840
rect 65 770 75 840
rect 35 725 75 770
rect 140 840 180 850
rect 140 770 150 840
rect 170 770 180 840
rect 140 760 180 770
rect 205 840 245 850
rect 205 770 215 840
rect 235 770 245 840
rect 205 740 245 770
rect 285 840 360 850
rect 285 770 295 840
rect 350 770 360 840
rect 285 760 360 770
rect 400 840 440 850
rect 400 770 410 840
rect 430 770 440 840
rect 35 705 45 725
rect 65 705 75 725
rect 35 695 75 705
rect 115 730 245 740
rect 115 710 215 730
rect 235 710 245 730
rect 400 740 440 770
rect 465 840 505 850
rect 465 770 475 840
rect 495 770 505 840
rect 465 760 505 770
rect 570 840 610 850
rect 570 770 580 840
rect 600 770 610 840
rect 400 730 445 740
rect 115 700 245 710
rect 275 705 365 715
rect -45 620 -5 630
rect -45 550 -35 620
rect -15 550 -5 620
rect -45 520 -5 550
rect 35 620 75 630
rect 35 550 45 620
rect 65 550 75 620
rect 35 540 75 550
rect 115 620 155 700
rect 275 680 285 705
rect 355 680 365 705
rect 400 710 410 730
rect 430 710 445 730
rect 400 700 445 710
rect 275 670 365 680
rect 115 550 125 620
rect 145 550 155 620
rect 115 520 155 550
rect -45 500 155 520
rect 180 620 220 630
rect 180 550 190 620
rect 210 550 220 620
rect 180 520 220 550
rect 260 620 300 630
rect 260 550 270 620
rect 290 550 300 620
rect 260 540 300 550
rect 340 620 380 630
rect 340 550 350 620
rect 370 550 380 620
rect 340 520 380 550
rect 180 500 380 520
rect 405 620 445 700
rect 570 725 610 770
rect 570 705 580 725
rect 600 705 610 725
rect 570 695 610 705
rect 405 550 415 620
rect 435 550 445 620
rect 405 520 445 550
rect 485 620 525 630
rect 485 550 495 620
rect 515 550 525 620
rect 485 540 525 550
rect 565 620 605 630
rect 565 550 575 620
rect 595 550 605 620
rect 565 520 605 550
rect 405 500 605 520
rect 135 470 175 480
rect 135 460 145 470
rect -135 450 145 460
rect 165 450 175 470
rect -135 440 175 450
rect 360 430 400 440
rect 360 420 370 430
rect -135 410 370 420
rect 390 410 400 430
rect -135 400 400 410
rect 520 390 560 400
rect 520 380 530 390
rect -135 370 530 380
rect 550 370 560 390
rect -135 360 560 370
rect -135 325 500 335
rect -135 315 470 325
rect 460 305 470 315
rect 490 305 500 325
rect 460 295 500 305
rect -135 285 40 295
rect -135 265 10 285
rect 30 265 40 285
rect -135 255 40 265
rect -135 225 145 235
rect -135 215 115 225
rect 105 205 115 215
rect 135 205 145 225
rect 105 195 145 205
rect 260 185 465 195
rect 260 165 270 185
rect 290 175 465 185
rect 290 165 300 175
rect -45 150 -5 160
rect -45 130 -35 150
rect -15 130 -5 150
rect -45 85 -5 130
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 -50 -5 15
rect 20 150 75 160
rect 260 155 300 165
rect 20 130 45 150
rect 65 130 75 150
rect 325 145 365 155
rect 325 135 335 145
rect 20 120 75 130
rect 150 125 335 135
rect 355 125 365 145
rect 20 85 60 120
rect 150 115 365 125
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect 85 -15 125 15
rect 150 85 190 115
rect 150 15 160 85
rect 180 15 190 85
rect 150 5 190 15
rect 215 85 255 95
rect 215 15 225 85
rect 245 15 255 85
rect 215 -15 255 15
rect 280 85 320 95
rect 280 15 290 85
rect 310 15 320 85
rect 280 5 320 15
rect 345 85 385 95
rect 345 15 355 85
rect 375 15 385 85
rect 85 -35 255 -15
rect 345 -15 385 15
rect 425 85 465 175
rect 570 150 610 160
rect 570 130 580 150
rect 600 130 610 150
rect 425 15 435 85
rect 455 15 465 85
rect 425 5 465 15
rect 505 85 545 95
rect 505 15 515 85
rect 535 15 545 85
rect 505 -15 545 15
rect 570 85 610 130
rect 570 15 580 85
rect 600 15 610 85
rect 570 5 610 15
rect 345 -35 545 -15
rect -45 -70 -35 -50
rect -15 -70 -5 -50
rect -45 -80 -5 -70
<< viali >>
rect -100 770 -80 840
rect -35 705 -15 725
rect 150 770 170 840
rect 295 770 350 840
rect 45 705 65 725
rect 475 770 495 840
rect 45 550 65 620
rect 285 680 355 705
rect 270 550 290 620
rect 580 705 600 725
rect 495 550 515 620
rect -35 130 -15 150
rect 45 130 65 150
rect 290 15 310 85
rect 580 130 600 150
<< metal1 >>
rect -135 840 685 855
rect -135 770 -100 840
rect -80 770 150 840
rect 170 770 295 840
rect 350 770 475 840
rect 495 770 685 840
rect -135 755 685 770
rect -135 500 -85 755
rect -50 735 0 740
rect -50 695 -45 735
rect -5 695 0 735
rect -50 690 0 695
rect 30 735 80 740
rect 30 695 35 735
rect 75 695 80 735
rect 565 735 615 740
rect 30 690 80 695
rect 270 705 370 720
rect 270 680 285 705
rect 355 680 370 705
rect 565 695 570 735
rect 610 695 615 735
rect 565 690 615 695
rect 270 635 370 680
rect -50 620 610 635
rect -50 550 45 620
rect 65 550 270 620
rect 290 550 495 620
rect 515 550 610 620
rect -50 535 610 550
rect -50 160 0 165
rect -50 120 -45 160
rect -5 120 0 160
rect -50 115 0 120
rect 30 160 80 165
rect 30 120 35 160
rect 75 120 80 160
rect 30 115 80 120
rect 270 100 370 535
rect 635 505 685 755
rect 565 160 615 165
rect 565 120 570 160
rect 610 120 615 160
rect 565 115 615 120
rect -135 85 685 100
rect -135 15 290 85
rect 310 15 685 85
rect -135 0 685 15
<< via1 >>
rect -45 725 -5 735
rect -45 705 -35 725
rect -35 705 -15 725
rect -15 705 -5 725
rect -45 695 -5 705
rect 35 725 75 735
rect 35 705 45 725
rect 45 705 65 725
rect 65 705 75 725
rect 35 695 75 705
rect 570 725 610 735
rect 570 705 580 725
rect 580 705 600 725
rect 600 705 610 725
rect 570 695 610 705
rect -45 150 -5 160
rect -45 130 -35 150
rect -35 130 -15 150
rect -15 130 -5 150
rect -45 120 -5 130
rect 35 150 75 160
rect 35 130 45 150
rect 45 130 65 150
rect 65 130 75 150
rect 35 120 75 130
rect 570 150 610 160
rect 570 130 580 150
rect 580 130 600 150
rect 600 130 610 150
rect 570 120 610 130
<< metal2 >>
rect -50 735 0 740
rect -50 695 -45 735
rect -5 695 0 735
rect -50 160 0 695
rect -50 120 -45 160
rect -5 120 0 160
rect -50 115 0 120
rect 30 735 80 740
rect 30 695 35 735
rect 75 695 80 735
rect 30 160 80 695
rect 30 120 35 160
rect 75 120 80 160
rect 30 115 80 120
rect 565 735 615 740
rect 565 695 570 735
rect 610 695 615 735
rect 565 160 615 695
rect 565 120 570 160
rect 610 120 615 160
rect 565 115 615 120
<< labels >>
flabel metal1 -135 50 -135 50 0 FreeSans 400 0 0 0 VN
port 2 nsew
flabel metal1 -135 550 -135 550 0 FreeSans 400 0 0 0 VP
port 3 nsew
flabel locali -135 225 -135 225 0 FreeSans 160 0 0 0 RST
port 4 nsew
flabel locali -135 275 -135 275 0 FreeSans 160 0 0 0 ENAD_n
port 5 nsew
flabel locali -135 325 -135 325 0 FreeSans 160 0 0 0 ENAD_p
port 6 nsew
flabel locali -135 450 -135 450 0 FreeSans 160 0 0 0 Ain
port 7 nsew
flabel locali -135 410 -135 410 0 FreeSans 160 0 0 0 Ui
port 8 nsew
flabel locali -135 370 -135 370 0 FreeSans 160 0 0 0 Vb
port 9 nsew
<< end >>
