magic
tech sky130A
timestamp 1702605448
<< nwell >>
rect -130 225 380 365
rect 270 195 380 225
rect 275 -50 380 195
<< nmos >>
rect -60 -25 -45 75
rect 5 -25 20 75
rect 170 -25 185 75
rect -60 -250 -45 -150
rect 5 -250 20 -150
rect 45 -250 60 -150
rect 110 -250 125 -150
rect 150 -250 165 -150
rect 215 -250 230 -150
<< pmos >>
rect -60 245 -45 345
rect 5 245 20 345
rect 45 245 60 345
rect 190 245 205 345
rect 230 245 245 345
rect 295 245 310 345
<< ndiff >>
rect -110 60 -60 75
rect -110 -10 -95 60
rect -75 -10 -60 60
rect -110 -25 -60 -10
rect -45 60 5 75
rect -45 -10 -30 60
rect -10 -10 5 60
rect -45 -25 5 -10
rect 20 60 70 75
rect 120 60 170 75
rect 20 -10 35 60
rect 55 -10 70 60
rect 120 -10 135 60
rect 155 -10 170 60
rect 20 -25 70 -10
rect 120 -25 170 -10
rect 185 60 235 75
rect 185 -10 200 60
rect 220 -10 235 60
rect 185 -25 235 -10
rect -110 -165 -60 -150
rect -110 -235 -95 -165
rect -75 -235 -60 -165
rect -110 -250 -60 -235
rect -45 -165 5 -150
rect -45 -235 -30 -165
rect -10 -235 5 -165
rect -45 -250 5 -235
rect 20 -250 45 -150
rect 60 -165 110 -150
rect 60 -235 75 -165
rect 95 -235 110 -165
rect 60 -250 110 -235
rect 125 -250 150 -150
rect 165 -165 215 -150
rect 165 -235 180 -165
rect 200 -235 215 -165
rect 165 -250 215 -235
rect 230 -165 280 -150
rect 230 -235 245 -165
rect 265 -235 280 -165
rect 230 -250 280 -235
<< pdiff >>
rect -110 330 -60 345
rect -110 260 -95 330
rect -75 260 -60 330
rect -110 245 -60 260
rect -45 330 5 345
rect -45 260 -30 330
rect -10 260 5 330
rect -45 245 5 260
rect 20 245 45 345
rect 60 330 110 345
rect 60 260 75 330
rect 95 260 110 330
rect 60 245 110 260
rect 140 330 190 345
rect 140 260 155 330
rect 175 260 190 330
rect 140 245 190 260
rect 205 245 230 345
rect 245 330 295 345
rect 245 260 260 330
rect 280 260 295 330
rect 245 245 295 260
rect 310 330 360 345
rect 310 260 325 330
rect 345 260 360 330
rect 310 245 360 260
<< ndiffc >>
rect -95 -10 -75 60
rect -30 -10 -10 60
rect 35 -10 55 60
rect 135 -10 155 60
rect 200 -10 220 60
rect -95 -235 -75 -165
rect -30 -235 -10 -165
rect 75 -235 95 -165
rect 180 -235 200 -165
rect 245 -235 265 -165
<< pdiffc >>
rect -95 260 -75 330
rect -30 260 -10 330
rect 75 260 95 330
rect 155 260 175 330
rect 260 260 280 330
rect 325 260 345 330
<< psubdiff >>
rect 70 60 120 75
rect 70 -10 90 60
rect 110 -10 120 60
rect 70 -25 120 -10
<< nsubdiff >>
rect 295 60 345 75
rect 295 -10 310 60
rect 330 -10 345 60
rect 295 -25 345 -10
<< psubdiffcont >>
rect 90 -10 110 60
<< nsubdiffcont >>
rect 310 -10 330 60
<< poly >>
rect 95 390 135 395
rect 95 370 105 390
rect 125 370 135 390
rect -60 345 -45 360
rect 5 345 20 360
rect 45 355 205 370
rect 45 345 60 355
rect 190 345 205 355
rect 230 345 245 360
rect 295 345 310 360
rect -60 235 -45 245
rect 5 235 20 245
rect -60 220 20 235
rect 45 230 60 245
rect 190 230 205 245
rect 230 235 245 245
rect 295 235 310 245
rect 230 220 310 235
rect -60 200 -50 220
rect -30 200 -20 220
rect -60 195 -20 200
rect 270 200 280 220
rect 300 200 310 220
rect 270 195 310 200
rect -130 185 -100 195
rect -130 165 -125 185
rect -105 170 -100 185
rect -105 165 185 170
rect -130 155 185 165
rect -130 115 -100 125
rect -130 95 -125 115
rect -105 100 -100 115
rect 80 120 120 125
rect 80 100 90 120
rect 110 100 120 120
rect -105 95 -45 100
rect -130 85 -45 95
rect -60 75 -45 85
rect 5 85 120 100
rect 5 75 20 85
rect 170 75 185 155
rect -60 -40 -45 -25
rect 5 -40 20 -25
rect 170 -40 185 -25
rect -115 -50 -85 -40
rect -115 -70 -110 -50
rect -90 -65 -85 -50
rect -90 -70 230 -65
rect -115 -80 230 -70
rect -85 -110 -45 -105
rect -85 -130 -75 -110
rect -55 -130 -45 -110
rect -85 -135 -45 -130
rect -60 -150 -45 -135
rect 5 -150 20 -135
rect 45 -150 60 -135
rect 110 -150 125 -135
rect 150 -150 165 -135
rect 215 -150 230 -80
rect -60 -265 -45 -250
rect 5 -315 20 -250
rect 45 -260 60 -250
rect 110 -260 125 -250
rect 45 -270 125 -260
rect 45 -275 75 -270
rect 65 -290 75 -275
rect 95 -275 125 -270
rect 95 -290 105 -275
rect 65 -295 105 -290
rect -20 -320 20 -315
rect -20 -340 -10 -320
rect 10 -340 20 -320
rect -20 -345 20 -340
rect 150 -315 165 -250
rect 215 -265 230 -250
rect 150 -320 190 -315
rect 150 -340 160 -320
rect 180 -340 190 -320
rect 150 -345 190 -340
<< polycont >>
rect 105 370 125 390
rect -50 200 -30 220
rect 280 200 300 220
rect -125 165 -105 185
rect -125 95 -105 115
rect 90 100 110 120
rect -110 -70 -90 -50
rect -75 -130 -55 -110
rect 75 -290 95 -270
rect -10 -340 10 -320
rect 160 -340 180 -320
<< locali >>
rect 95 390 135 395
rect -130 370 105 390
rect 125 370 135 390
rect 95 365 135 370
rect -105 330 -60 340
rect -105 260 -95 330
rect -75 260 -60 330
rect -105 250 -60 260
rect -40 330 0 340
rect -40 260 -30 330
rect -10 260 0 330
rect -40 250 0 260
rect 65 330 105 340
rect 65 260 75 330
rect 95 260 105 330
rect -80 225 -60 250
rect 65 225 105 260
rect -80 220 -20 225
rect -80 200 -50 220
rect -30 200 -20 220
rect 65 205 75 225
rect 95 205 105 225
rect 65 200 105 205
rect 145 330 185 340
rect 145 260 155 330
rect 175 260 185 330
rect 145 225 185 260
rect 250 330 290 340
rect 250 260 260 330
rect 280 260 290 330
rect 250 250 290 260
rect 315 330 355 340
rect 315 260 325 330
rect 345 260 355 330
rect 315 250 355 260
rect 325 225 345 250
rect 145 205 155 225
rect 175 205 185 225
rect 145 200 185 205
rect 270 220 345 225
rect 270 200 280 220
rect 300 200 345 220
rect -80 195 -20 200
rect 270 195 345 200
rect -130 185 -100 195
rect -130 165 -125 185
rect -105 165 -100 185
rect -130 155 -100 165
rect -130 115 -100 125
rect -130 95 -125 115
rect -105 95 -100 115
rect -130 85 -100 95
rect -80 65 -60 195
rect 270 180 290 195
rect 35 160 290 180
rect 35 70 55 160
rect 80 120 380 125
rect 80 100 90 120
rect 110 100 380 120
rect 80 95 380 100
rect -105 60 -60 65
rect -105 -10 -95 60
rect -75 -10 -60 60
rect -105 -20 -60 -10
rect -40 60 0 70
rect -40 -10 -30 60
rect -10 -10 0 60
rect -40 -20 0 -10
rect 25 60 65 70
rect 25 -10 35 60
rect 55 -10 65 60
rect 25 -20 65 -10
rect 85 60 165 70
rect 85 -10 90 60
rect 110 -10 135 60
rect 155 -10 165 60
rect 85 -20 165 -10
rect 190 60 230 70
rect 190 -10 200 60
rect 220 -10 230 60
rect 190 -20 230 -10
rect 300 60 340 70
rect 300 -10 310 60
rect 330 -10 340 60
rect 300 -20 340 -10
rect -30 -40 -10 -20
rect 200 -40 220 -20
rect -130 -50 -85 -40
rect -130 -70 -110 -50
rect -90 -70 -85 -50
rect -30 -60 220 -40
rect -130 -80 -85 -70
rect -25 -95 5 -85
rect -130 -110 -45 -105
rect -130 -130 -75 -110
rect -55 -130 -45 -110
rect -130 -135 -45 -130
rect -25 -115 -20 -95
rect 0 -115 5 -95
rect -25 -125 5 -115
rect 165 -100 195 -90
rect 165 -120 170 -100
rect 190 -120 195 -100
rect -25 -155 0 -125
rect 165 -130 195 -120
rect 170 -155 195 -130
rect -105 -165 -65 -155
rect -105 -235 -95 -165
rect -75 -235 -65 -165
rect -105 -265 -65 -235
rect -40 -165 0 -155
rect -40 -235 -30 -165
rect -10 -235 0 -165
rect -40 -245 0 -235
rect 65 -165 105 -155
rect 65 -235 75 -165
rect 95 -235 105 -165
rect 65 -245 105 -235
rect 170 -165 210 -155
rect 170 -235 180 -165
rect 200 -235 210 -165
rect 170 -245 210 -235
rect 235 -165 275 -155
rect 235 -235 245 -165
rect 265 -235 275 -165
rect 235 -265 275 -235
rect -105 -270 275 -265
rect -105 -290 75 -270
rect 95 -290 275 -270
rect -105 -295 275 -290
rect -130 -320 380 -315
rect -130 -340 -10 -320
rect 10 -340 160 -320
rect 180 -340 380 -320
rect -130 -345 380 -340
<< viali >>
rect -30 260 -10 330
rect 75 205 95 225
rect 260 260 280 330
rect 155 205 175 225
rect 90 -10 110 60
rect 135 -10 155 60
rect 310 -10 330 60
rect -20 -115 0 -95
rect 170 -120 190 -100
rect 75 -235 95 -165
<< metal1 >>
rect -130 330 380 340
rect -130 260 -30 330
rect -10 260 260 330
rect 280 260 380 330
rect -130 250 380 260
rect -25 225 105 230
rect -25 205 75 225
rect 95 205 105 225
rect -25 200 105 205
rect 145 225 225 230
rect 145 205 155 225
rect 175 205 225 225
rect 145 200 225 205
rect -25 -95 5 200
rect -25 -115 -20 -95
rect 0 -115 5 -95
rect -25 -125 5 -115
rect 85 60 165 70
rect 85 -10 90 60
rect 110 -10 135 60
rect 155 -10 165 60
rect 85 -20 165 -10
rect 85 -155 135 -20
rect 195 -90 225 200
rect 300 60 340 250
rect 300 -10 310 60
rect 330 -10 340 60
rect 300 -20 340 -10
rect 165 -100 225 -90
rect 165 -120 170 -100
rect 190 -120 225 -100
rect 165 -130 225 -120
rect -130 -165 380 -155
rect -130 -235 75 -165
rect 95 -235 380 -165
rect -130 -245 380 -235
<< labels >>
rlabel locali -130 -60 -130 -60 7 Vinv_n
port 5 w
rlabel locali -130 -120 -130 -120 7 Vinv_p
port 6 w
rlabel metal1 -130 -200 -130 -200 7 VN
port 7 w
rlabel locali -130 -330 -130 -330 7 Vcn
port 8 w
rlabel locali -130 380 -130 380 7 Vcp
port 1 w
rlabel metal1 -130 295 -130 295 7 VP
port 2 w
rlabel locali -130 175 -130 175 7 Vb
port 3 w
rlabel locali -130 105 -130 105 7 Vin_n
port 4 w
rlabel locali 380 110 380 110 3 Vin_p
port 9 e
<< end >>
