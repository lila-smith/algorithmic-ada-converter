magic
tech sky130A
timestamp 1702706444
<< nwell >>
rect -135 715 620 855
<< nmos >>
rect 95 535 110 635
rect 160 535 175 635
rect 225 535 240 635
rect 395 535 410 635
rect 460 535 475 635
rect 0 0 15 100
rect 65 0 80 100
rect 130 0 145 100
rect 195 0 210 100
rect 260 0 275 100
rect 325 0 340 100
rect 390 0 405 100
rect 535 0 550 100
<< pmos >>
rect -65 735 -50 835
rect 80 735 95 835
rect 120 735 135 835
rect 185 735 200 835
rect 430 735 445 835
rect 495 735 510 835
rect 535 735 550 835
<< ndiff >>
rect 45 620 95 635
rect 45 550 60 620
rect 80 550 95 620
rect 45 535 95 550
rect 110 620 160 635
rect 110 550 125 620
rect 145 550 160 620
rect 110 535 160 550
rect 175 620 225 635
rect 175 550 190 620
rect 210 550 225 620
rect 175 535 225 550
rect 240 620 290 635
rect 345 620 395 635
rect 240 550 255 620
rect 280 550 290 620
rect 345 550 360 620
rect 380 550 395 620
rect 240 535 290 550
rect 345 535 395 550
rect 410 620 460 635
rect 410 550 425 620
rect 445 550 460 620
rect 410 535 460 550
rect 475 620 525 635
rect 475 550 490 620
rect 510 550 525 620
rect 475 535 525 550
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 145 85 195 100
rect 145 15 160 85
rect 180 15 195 85
rect 145 0 195 15
rect 210 85 260 100
rect 210 15 225 85
rect 245 15 260 85
rect 210 0 260 15
rect 275 85 325 100
rect 275 15 290 85
rect 310 15 325 85
rect 275 0 325 15
rect 340 85 390 100
rect 340 15 355 85
rect 375 15 390 85
rect 340 0 390 15
rect 405 85 455 100
rect 405 15 420 85
rect 440 15 455 85
rect 405 0 455 15
rect 485 85 535 100
rect 485 15 500 85
rect 520 15 535 85
rect 485 0 535 15
rect 550 85 600 100
rect 550 15 565 85
rect 585 15 600 85
rect 550 0 600 15
<< pdiff >>
rect -115 820 -65 835
rect -115 750 -100 820
rect -80 750 -65 820
rect -115 735 -65 750
rect -50 820 0 835
rect -50 750 -35 820
rect -15 750 0 820
rect -50 735 0 750
rect 30 820 80 835
rect 30 750 45 820
rect 65 750 80 820
rect 30 735 80 750
rect 95 735 120 835
rect 135 820 185 835
rect 135 750 150 820
rect 170 750 185 820
rect 135 735 185 750
rect 200 820 250 835
rect 200 750 215 820
rect 235 750 250 820
rect 200 735 250 750
rect 380 820 430 835
rect 380 750 395 820
rect 415 750 430 820
rect 380 735 430 750
rect 445 820 495 835
rect 445 750 460 820
rect 480 750 495 820
rect 445 735 495 750
rect 510 735 535 835
rect 550 820 600 835
rect 550 750 565 820
rect 585 750 600 820
rect 550 735 600 750
<< ndiffc >>
rect 60 550 80 620
rect 125 550 145 620
rect 190 550 210 620
rect 255 550 280 620
rect 360 550 380 620
rect 425 550 445 620
rect 490 550 510 620
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
rect 160 15 180 85
rect 225 15 245 85
rect 290 15 310 85
rect 355 15 375 85
rect 420 15 440 85
rect 500 15 520 85
rect 565 15 585 85
<< pdiffc >>
rect -100 750 -80 820
rect -35 750 -15 820
rect 45 750 65 820
rect 150 750 170 820
rect 215 750 235 820
rect 395 750 415 820
rect 460 750 480 820
rect 565 750 585 820
<< psubdiff >>
rect 290 620 345 635
rect 290 550 300 620
rect 325 550 345 620
rect 290 535 345 550
<< nsubdiff >>
rect 280 820 350 835
rect 280 750 295 820
rect 335 750 350 820
rect 280 735 350 750
<< psubdiffcont >>
rect 300 550 325 620
<< nsubdiffcont >>
rect 295 750 335 820
<< poly >>
rect 55 880 550 890
rect 55 860 65 880
rect 85 875 550 880
rect 85 860 95 875
rect 55 850 95 860
rect -65 835 -50 850
rect 80 835 95 850
rect 120 835 135 850
rect 185 835 200 850
rect 430 835 445 850
rect 495 835 510 850
rect 535 835 550 875
rect -65 715 -50 735
rect 80 720 95 735
rect 120 720 135 735
rect 185 720 200 735
rect 430 720 445 735
rect 495 720 510 735
rect 535 720 550 735
rect -75 700 -50 715
rect 120 710 245 720
rect 120 705 215 710
rect -75 295 -60 700
rect 205 690 215 705
rect 235 690 245 710
rect 205 680 245 690
rect 385 710 510 720
rect 385 690 395 710
rect 415 705 510 710
rect 415 690 425 705
rect 385 680 425 690
rect 95 635 110 650
rect 160 635 175 650
rect 225 635 240 650
rect 395 635 410 650
rect 460 635 475 650
rect 95 375 110 535
rect 160 480 175 535
rect 135 470 175 480
rect 135 450 145 470
rect 165 450 175 470
rect 135 440 175 450
rect 225 375 240 535
rect 395 440 410 535
rect 370 400 410 440
rect 460 400 475 535
rect 450 390 490 400
rect 450 375 460 390
rect 95 370 460 375
rect 480 370 490 390
rect 95 360 490 370
rect 460 325 500 335
rect 460 305 470 325
rect 490 305 500 325
rect 460 295 500 305
rect -75 285 210 295
rect -75 280 10 285
rect 0 265 10 280
rect 30 280 210 285
rect 30 265 40 280
rect 0 255 40 265
rect 0 100 15 255
rect 105 225 145 235
rect 105 205 115 225
rect 135 205 145 225
rect 105 195 145 205
rect 65 100 80 115
rect 130 100 145 195
rect 195 100 210 280
rect 260 185 300 195
rect 260 165 270 185
rect 290 165 300 185
rect 260 155 300 165
rect 260 100 275 155
rect 325 145 365 155
rect 325 125 335 145
rect 355 125 365 145
rect 460 125 475 295
rect 325 115 365 125
rect 325 100 340 115
rect 390 110 475 125
rect 390 100 405 110
rect 535 100 550 115
rect 0 -15 15 0
rect 65 -40 80 0
rect 130 -15 145 0
rect 195 -15 210 0
rect 260 -15 275 0
rect 325 -15 340 0
rect 390 -15 405 0
rect 535 -40 550 0
rect -45 -50 550 -40
rect -45 -70 -35 -50
rect -15 -55 550 -50
rect -15 -70 -5 -55
rect -45 -80 -5 -70
<< polycont >>
rect 65 860 85 880
rect 215 690 235 710
rect 395 690 415 710
rect 145 450 165 470
rect 460 370 480 390
rect 470 305 490 325
rect 10 265 30 285
rect 115 205 135 225
rect 270 165 290 185
rect 335 125 355 145
rect -35 -70 -15 -50
<< locali >>
rect -135 880 95 890
rect -135 870 65 880
rect 55 860 65 870
rect 85 860 95 880
rect 55 850 95 860
rect -110 820 -70 830
rect -110 750 -100 820
rect -80 750 -70 820
rect -110 740 -70 750
rect -45 820 -5 830
rect -45 750 -35 820
rect -15 750 -5 820
rect -45 720 -5 750
rect -70 710 -5 720
rect -70 690 -60 710
rect -40 690 -5 710
rect -70 680 -5 690
rect 35 820 75 830
rect 35 750 45 820
rect 65 750 75 820
rect 35 710 75 750
rect 140 820 180 830
rect 140 750 150 820
rect 170 750 180 820
rect 140 740 180 750
rect 205 820 245 830
rect 205 750 215 820
rect 235 750 245 820
rect 205 720 245 750
rect 285 820 345 830
rect 285 750 295 820
rect 335 750 345 820
rect 285 740 345 750
rect 385 820 425 830
rect 385 750 395 820
rect 415 750 425 820
rect 35 690 45 710
rect 65 690 75 710
rect 35 680 75 690
rect 115 710 245 720
rect 115 690 215 710
rect 235 690 245 710
rect 115 680 245 690
rect 385 720 425 750
rect 450 820 490 830
rect 450 750 460 820
rect 480 750 490 820
rect 450 740 490 750
rect 555 820 595 830
rect 555 750 565 820
rect 585 750 595 820
rect 385 710 455 720
rect 385 690 395 710
rect 415 690 455 710
rect 385 680 455 690
rect 555 710 595 750
rect 555 690 565 710
rect 585 690 595 710
rect 555 680 595 690
rect 50 620 90 630
rect 50 550 60 620
rect 80 550 90 620
rect 50 540 90 550
rect 115 620 155 680
rect 115 550 125 620
rect 145 550 155 620
rect 115 540 155 550
rect 180 620 220 630
rect 180 550 190 620
rect 210 550 220 620
rect 180 520 220 550
rect 245 620 330 630
rect 245 550 255 620
rect 280 550 300 620
rect 325 550 330 620
rect 245 540 330 550
rect 350 620 390 630
rect 350 550 360 620
rect 380 550 390 620
rect 350 520 390 550
rect 415 620 455 680
rect 415 550 425 620
rect 445 550 455 620
rect 415 540 455 550
rect 480 620 520 630
rect 480 550 490 620
rect 510 550 520 620
rect 480 540 520 550
rect 180 500 390 520
rect 135 470 175 480
rect 135 460 145 470
rect -135 450 145 460
rect 165 450 175 470
rect -135 440 175 450
rect 370 420 410 440
rect -135 400 410 420
rect 450 390 490 400
rect 450 380 460 390
rect -135 370 460 380
rect 480 370 490 390
rect -135 360 490 370
rect -135 325 500 335
rect -135 315 470 325
rect 460 305 470 315
rect 490 305 500 325
rect 460 295 500 305
rect -135 285 40 295
rect -135 265 10 285
rect 30 265 40 285
rect -135 255 40 265
rect -135 225 145 235
rect -135 215 115 225
rect 105 205 115 215
rect 135 205 145 225
rect 105 195 145 205
rect 260 185 450 195
rect 260 175 270 185
rect 150 165 270 175
rect 290 175 450 185
rect 290 165 300 175
rect 150 155 300 165
rect -70 145 -5 155
rect -70 125 -60 145
rect -40 125 -5 145
rect -70 115 -5 125
rect -45 85 -5 115
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 -50 -5 15
rect 20 145 60 155
rect 20 125 30 145
rect 50 125 60 145
rect 20 85 60 125
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect 85 -15 125 15
rect 150 85 190 155
rect 325 145 365 155
rect 325 135 335 145
rect 150 15 160 85
rect 180 15 190 85
rect 150 5 190 15
rect 215 125 335 135
rect 355 125 365 145
rect 215 115 365 125
rect 215 95 250 115
rect 215 85 255 95
rect 215 15 225 85
rect 245 15 255 85
rect 215 -15 255 15
rect 280 85 320 95
rect 280 15 290 85
rect 310 15 320 85
rect 280 5 320 15
rect 345 85 385 95
rect 345 15 355 85
rect 375 15 385 85
rect 85 -35 255 -15
rect 345 -15 385 15
rect 410 85 450 175
rect 555 145 595 155
rect 555 125 565 145
rect 585 125 595 145
rect 410 15 420 85
rect 440 15 450 85
rect 410 5 450 15
rect 490 85 530 95
rect 490 15 500 85
rect 520 15 530 85
rect 490 -15 530 15
rect 555 85 595 125
rect 555 15 565 85
rect 585 15 595 85
rect 555 5 595 15
rect 345 -35 530 -15
rect -45 -70 -35 -50
rect -15 -70 -5 -50
rect -45 -80 -5 -70
<< viali >>
rect -100 750 -80 820
rect -60 690 -40 710
rect 150 750 170 820
rect 295 750 335 820
rect 45 690 65 710
rect 460 750 480 820
rect 565 690 585 710
rect 60 550 80 620
rect 255 550 280 620
rect 300 550 325 620
rect 490 550 510 620
rect -60 125 -40 145
rect 30 125 50 145
rect 290 15 310 85
rect 565 125 585 145
<< metal1 >>
rect -135 820 670 835
rect -135 750 -100 820
rect -80 750 150 820
rect 170 750 295 820
rect 335 750 460 820
rect 480 750 670 820
rect -135 735 670 750
rect -135 500 -85 735
rect -70 710 -30 720
rect -70 690 -60 710
rect -40 690 -30 710
rect -70 145 -30 690
rect -70 125 -60 145
rect -40 125 -30 145
rect -70 115 -30 125
rect -15 710 75 720
rect -15 690 45 710
rect 65 690 75 710
rect -15 680 75 690
rect 555 710 595 720
rect 555 690 565 710
rect 585 690 595 710
rect -15 155 25 680
rect 45 620 525 635
rect 45 550 60 620
rect 80 550 255 620
rect 280 550 300 620
rect 325 550 490 620
rect 510 550 525 620
rect 45 535 525 550
rect -15 145 60 155
rect -15 125 30 145
rect 50 125 60 145
rect -15 115 60 125
rect 270 100 370 535
rect 555 145 595 690
rect 620 500 670 735
rect 555 125 565 145
rect 585 125 595 145
rect 555 115 595 125
rect -135 85 670 100
rect -135 15 290 85
rect 310 15 670 85
rect -135 0 670 15
<< labels >>
flabel metal1 -135 50 -135 50 0 FreeSans 400 0 0 0 VN
port 2 nsew
flabel metal1 -135 550 -135 550 0 FreeSans 400 0 0 0 VP
port 3 nsew
flabel locali -135 225 -135 225 0 FreeSans 160 0 0 0 RST
port 4 nsew
flabel locali -135 275 -135 275 0 FreeSans 160 0 0 0 ENAD_n
port 5 nsew
flabel locali -135 325 -135 325 0 FreeSans 160 0 0 0 ENAD_p
port 6 nsew
flabel locali -135 450 -135 450 0 FreeSans 160 0 0 0 Ain
port 7 nsew
flabel locali -135 410 -135 410 0 FreeSans 160 0 0 0 Ui
port 8 nsew
flabel locali -135 370 -135 370 0 FreeSans 160 0 0 0 Vb
port 9 nsew
<< end >>
